TITRE
░
Corp\n
du text
░
imageType.png
░
lienExemple
ExempleLien